`default_nettype none

module abus_rr #(

) (

);

endmodule