
localparam [1:0] S_IDLE  = 2'b00;
localparam [1:0] S_WRITE = 2'b01;
localparam [1:0] S_READ  = 2'b10;
localparam [1:0] S_ABORT = 2'b11;
