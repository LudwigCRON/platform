localparam NONE_ADR =   0;
localparam RO1_ADR  =   1;
localparam RO2_ADR  =   2;
localparam RW1_ADR  =   4;
localparam RW2_ADR  =   8;
localparam RW3_ADR  =  16;
localparam RWE1_ADR =  32;
localparam RWE2_ADR =  64;
localparam RWE3_ADR = 128;
localparam WO1_ADR  = 256;
localparam MIX1_ADR = 512;
localparam MIX2_ADR =1024;