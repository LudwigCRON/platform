
localparam [1:0] S_IDLE   = 2'b00;
localparam [1:0] S_WAIT   = 2'b01;
localparam [1:0] S_SAMPLE = 2'b11;